VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_example
  CLASS BLOCK ;
  FOREIGN user_proj_example ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 3000.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 99.320 200.000 99.920 ;
    END
  END io_in[0]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 699.080 200.000 699.680 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 1298.840 200.000 1299.440 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 1898.600 200.000 1899.200 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 2498.360 200.000 2498.960 ;
    END
  END io_in[4]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 499.160 200.000 499.760 ;
    END
  END io_oeb[0]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 1098.920 200.000 1099.520 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 1698.680 200.000 1699.280 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 2298.440 200.000 2299.040 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 2898.200 200.000 2898.800 ;
    END
  END io_oeb[4]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 299.240 200.000 299.840 ;
    END
  END io_out[0]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 899.000 200.000 899.600 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 1498.760 200.000 1499.360 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 2098.520 200.000 2099.120 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 2698.280 200.000 2698.880 ;
    END
  END io_out[4]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 2986.800 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 2986.800 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 149.590 0.000 149.870 4.000 ;
    END
  END wb_rst_i
  OBS
      LAYER nwell ;
        RECT 5.330 2982.425 194.310 2985.255 ;
        RECT 5.330 2976.985 194.310 2979.815 ;
        RECT 5.330 2971.545 194.310 2974.375 ;
        RECT 5.330 2966.105 194.310 2968.935 ;
        RECT 5.330 2960.665 194.310 2963.495 ;
        RECT 5.330 2955.225 194.310 2958.055 ;
        RECT 5.330 2949.785 194.310 2952.615 ;
        RECT 5.330 2944.345 194.310 2947.175 ;
        RECT 5.330 2938.905 194.310 2941.735 ;
        RECT 5.330 2933.465 194.310 2936.295 ;
        RECT 5.330 2928.025 194.310 2930.855 ;
        RECT 5.330 2922.585 194.310 2925.415 ;
        RECT 5.330 2917.145 194.310 2919.975 ;
        RECT 5.330 2911.705 194.310 2914.535 ;
        RECT 5.330 2906.265 194.310 2909.095 ;
        RECT 5.330 2900.825 194.310 2903.655 ;
        RECT 5.330 2895.385 194.310 2898.215 ;
        RECT 5.330 2889.945 194.310 2892.775 ;
        RECT 5.330 2884.505 194.310 2887.335 ;
        RECT 5.330 2879.065 194.310 2881.895 ;
        RECT 5.330 2873.625 194.310 2876.455 ;
        RECT 5.330 2868.185 194.310 2871.015 ;
        RECT 5.330 2862.745 194.310 2865.575 ;
        RECT 5.330 2857.305 194.310 2860.135 ;
        RECT 5.330 2851.865 194.310 2854.695 ;
        RECT 5.330 2846.425 194.310 2849.255 ;
        RECT 5.330 2840.985 194.310 2843.815 ;
        RECT 5.330 2835.545 194.310 2838.375 ;
        RECT 5.330 2830.105 194.310 2832.935 ;
        RECT 5.330 2824.665 194.310 2827.495 ;
        RECT 5.330 2819.225 194.310 2822.055 ;
        RECT 5.330 2813.785 194.310 2816.615 ;
        RECT 5.330 2808.345 194.310 2811.175 ;
        RECT 5.330 2802.905 194.310 2805.735 ;
        RECT 5.330 2797.465 194.310 2800.295 ;
        RECT 5.330 2792.025 194.310 2794.855 ;
        RECT 5.330 2786.585 194.310 2789.415 ;
        RECT 5.330 2781.145 194.310 2783.975 ;
        RECT 5.330 2775.705 194.310 2778.535 ;
        RECT 5.330 2770.265 194.310 2773.095 ;
        RECT 5.330 2764.825 194.310 2767.655 ;
        RECT 5.330 2759.385 194.310 2762.215 ;
        RECT 5.330 2753.945 194.310 2756.775 ;
        RECT 5.330 2748.505 194.310 2751.335 ;
        RECT 5.330 2743.065 194.310 2745.895 ;
        RECT 5.330 2737.625 194.310 2740.455 ;
        RECT 5.330 2732.185 194.310 2735.015 ;
        RECT 5.330 2726.745 194.310 2729.575 ;
        RECT 5.330 2721.305 194.310 2724.135 ;
        RECT 5.330 2715.865 194.310 2718.695 ;
        RECT 5.330 2710.425 194.310 2713.255 ;
        RECT 5.330 2704.985 194.310 2707.815 ;
        RECT 5.330 2699.545 194.310 2702.375 ;
        RECT 5.330 2694.105 194.310 2696.935 ;
        RECT 5.330 2688.665 194.310 2691.495 ;
        RECT 5.330 2683.225 194.310 2686.055 ;
        RECT 5.330 2677.785 194.310 2680.615 ;
        RECT 5.330 2672.345 194.310 2675.175 ;
        RECT 5.330 2666.905 194.310 2669.735 ;
        RECT 5.330 2661.465 194.310 2664.295 ;
        RECT 5.330 2656.025 194.310 2658.855 ;
        RECT 5.330 2650.585 194.310 2653.415 ;
        RECT 5.330 2645.145 194.310 2647.975 ;
        RECT 5.330 2639.705 194.310 2642.535 ;
        RECT 5.330 2634.265 194.310 2637.095 ;
        RECT 5.330 2628.825 194.310 2631.655 ;
        RECT 5.330 2623.385 194.310 2626.215 ;
        RECT 5.330 2617.945 194.310 2620.775 ;
        RECT 5.330 2612.505 194.310 2615.335 ;
        RECT 5.330 2607.065 194.310 2609.895 ;
        RECT 5.330 2601.625 194.310 2604.455 ;
        RECT 5.330 2596.185 194.310 2599.015 ;
        RECT 5.330 2590.745 194.310 2593.575 ;
        RECT 5.330 2585.305 194.310 2588.135 ;
        RECT 5.330 2579.865 194.310 2582.695 ;
        RECT 5.330 2574.425 194.310 2577.255 ;
        RECT 5.330 2568.985 194.310 2571.815 ;
        RECT 5.330 2563.545 194.310 2566.375 ;
        RECT 5.330 2558.105 194.310 2560.935 ;
        RECT 5.330 2552.665 194.310 2555.495 ;
        RECT 5.330 2547.225 194.310 2550.055 ;
        RECT 5.330 2541.785 194.310 2544.615 ;
        RECT 5.330 2536.345 194.310 2539.175 ;
        RECT 5.330 2530.905 194.310 2533.735 ;
        RECT 5.330 2525.465 194.310 2528.295 ;
        RECT 5.330 2520.025 194.310 2522.855 ;
        RECT 5.330 2514.585 194.310 2517.415 ;
        RECT 5.330 2509.145 194.310 2511.975 ;
        RECT 5.330 2503.705 194.310 2506.535 ;
        RECT 5.330 2498.265 194.310 2501.095 ;
        RECT 5.330 2492.825 194.310 2495.655 ;
        RECT 5.330 2487.385 194.310 2490.215 ;
        RECT 5.330 2481.945 194.310 2484.775 ;
        RECT 5.330 2476.505 194.310 2479.335 ;
        RECT 5.330 2471.065 194.310 2473.895 ;
        RECT 5.330 2465.625 194.310 2468.455 ;
        RECT 5.330 2460.185 194.310 2463.015 ;
        RECT 5.330 2454.745 194.310 2457.575 ;
        RECT 5.330 2449.305 194.310 2452.135 ;
        RECT 5.330 2443.865 194.310 2446.695 ;
        RECT 5.330 2438.425 194.310 2441.255 ;
        RECT 5.330 2432.985 194.310 2435.815 ;
        RECT 5.330 2427.545 194.310 2430.375 ;
        RECT 5.330 2422.105 194.310 2424.935 ;
        RECT 5.330 2416.665 194.310 2419.495 ;
        RECT 5.330 2411.225 194.310 2414.055 ;
        RECT 5.330 2405.785 194.310 2408.615 ;
        RECT 5.330 2400.345 194.310 2403.175 ;
        RECT 5.330 2394.905 194.310 2397.735 ;
        RECT 5.330 2389.465 194.310 2392.295 ;
        RECT 5.330 2384.025 194.310 2386.855 ;
        RECT 5.330 2378.585 194.310 2381.415 ;
        RECT 5.330 2373.145 194.310 2375.975 ;
        RECT 5.330 2367.705 194.310 2370.535 ;
        RECT 5.330 2362.265 194.310 2365.095 ;
        RECT 5.330 2356.825 194.310 2359.655 ;
        RECT 5.330 2351.385 194.310 2354.215 ;
        RECT 5.330 2345.945 194.310 2348.775 ;
        RECT 5.330 2340.505 194.310 2343.335 ;
        RECT 5.330 2335.065 194.310 2337.895 ;
        RECT 5.330 2329.625 194.310 2332.455 ;
        RECT 5.330 2324.185 194.310 2327.015 ;
        RECT 5.330 2318.745 194.310 2321.575 ;
        RECT 5.330 2313.305 194.310 2316.135 ;
        RECT 5.330 2307.865 194.310 2310.695 ;
        RECT 5.330 2302.425 194.310 2305.255 ;
        RECT 5.330 2296.985 194.310 2299.815 ;
        RECT 5.330 2291.545 194.310 2294.375 ;
        RECT 5.330 2286.105 194.310 2288.935 ;
        RECT 5.330 2280.665 194.310 2283.495 ;
        RECT 5.330 2275.225 194.310 2278.055 ;
        RECT 5.330 2269.785 194.310 2272.615 ;
        RECT 5.330 2264.345 194.310 2267.175 ;
        RECT 5.330 2258.905 194.310 2261.735 ;
        RECT 5.330 2253.465 194.310 2256.295 ;
        RECT 5.330 2248.025 194.310 2250.855 ;
        RECT 5.330 2242.585 194.310 2245.415 ;
        RECT 5.330 2237.145 194.310 2239.975 ;
        RECT 5.330 2231.705 194.310 2234.535 ;
        RECT 5.330 2226.265 194.310 2229.095 ;
        RECT 5.330 2220.825 194.310 2223.655 ;
        RECT 5.330 2215.385 194.310 2218.215 ;
        RECT 5.330 2209.945 194.310 2212.775 ;
        RECT 5.330 2204.505 194.310 2207.335 ;
        RECT 5.330 2199.065 194.310 2201.895 ;
        RECT 5.330 2193.625 194.310 2196.455 ;
        RECT 5.330 2188.185 194.310 2191.015 ;
        RECT 5.330 2182.745 194.310 2185.575 ;
        RECT 5.330 2177.305 194.310 2180.135 ;
        RECT 5.330 2171.865 194.310 2174.695 ;
        RECT 5.330 2166.425 194.310 2169.255 ;
        RECT 5.330 2160.985 194.310 2163.815 ;
        RECT 5.330 2155.545 194.310 2158.375 ;
        RECT 5.330 2150.105 194.310 2152.935 ;
        RECT 5.330 2144.665 194.310 2147.495 ;
        RECT 5.330 2139.225 194.310 2142.055 ;
        RECT 5.330 2133.785 194.310 2136.615 ;
        RECT 5.330 2128.345 194.310 2131.175 ;
        RECT 5.330 2122.905 194.310 2125.735 ;
        RECT 5.330 2117.465 194.310 2120.295 ;
        RECT 5.330 2112.025 194.310 2114.855 ;
        RECT 5.330 2106.585 194.310 2109.415 ;
        RECT 5.330 2101.145 194.310 2103.975 ;
        RECT 5.330 2095.705 194.310 2098.535 ;
        RECT 5.330 2090.265 194.310 2093.095 ;
        RECT 5.330 2084.825 194.310 2087.655 ;
        RECT 5.330 2079.385 194.310 2082.215 ;
        RECT 5.330 2073.945 194.310 2076.775 ;
        RECT 5.330 2068.505 194.310 2071.335 ;
        RECT 5.330 2063.065 194.310 2065.895 ;
        RECT 5.330 2057.625 194.310 2060.455 ;
        RECT 5.330 2052.185 194.310 2055.015 ;
        RECT 5.330 2046.745 194.310 2049.575 ;
        RECT 5.330 2041.305 194.310 2044.135 ;
        RECT 5.330 2035.865 194.310 2038.695 ;
        RECT 5.330 2030.425 194.310 2033.255 ;
        RECT 5.330 2024.985 194.310 2027.815 ;
        RECT 5.330 2019.545 194.310 2022.375 ;
        RECT 5.330 2014.105 194.310 2016.935 ;
        RECT 5.330 2008.665 194.310 2011.495 ;
        RECT 5.330 2003.225 194.310 2006.055 ;
        RECT 5.330 1997.785 194.310 2000.615 ;
        RECT 5.330 1992.345 194.310 1995.175 ;
        RECT 5.330 1986.905 194.310 1989.735 ;
        RECT 5.330 1981.465 194.310 1984.295 ;
        RECT 5.330 1976.025 194.310 1978.855 ;
        RECT 5.330 1970.585 194.310 1973.415 ;
        RECT 5.330 1965.145 194.310 1967.975 ;
        RECT 5.330 1959.705 194.310 1962.535 ;
        RECT 5.330 1954.265 194.310 1957.095 ;
        RECT 5.330 1948.825 194.310 1951.655 ;
        RECT 5.330 1943.385 194.310 1946.215 ;
        RECT 5.330 1937.945 194.310 1940.775 ;
        RECT 5.330 1932.505 194.310 1935.335 ;
        RECT 5.330 1927.065 194.310 1929.895 ;
        RECT 5.330 1921.625 194.310 1924.455 ;
        RECT 5.330 1916.185 194.310 1919.015 ;
        RECT 5.330 1910.745 194.310 1913.575 ;
        RECT 5.330 1905.305 194.310 1908.135 ;
        RECT 5.330 1899.865 194.310 1902.695 ;
        RECT 5.330 1894.425 194.310 1897.255 ;
        RECT 5.330 1888.985 194.310 1891.815 ;
        RECT 5.330 1883.545 194.310 1886.375 ;
        RECT 5.330 1878.105 194.310 1880.935 ;
        RECT 5.330 1872.665 194.310 1875.495 ;
        RECT 5.330 1867.225 194.310 1870.055 ;
        RECT 5.330 1861.785 194.310 1864.615 ;
        RECT 5.330 1856.345 194.310 1859.175 ;
        RECT 5.330 1850.905 194.310 1853.735 ;
        RECT 5.330 1845.465 194.310 1848.295 ;
        RECT 5.330 1840.025 194.310 1842.855 ;
        RECT 5.330 1834.585 194.310 1837.415 ;
        RECT 5.330 1829.145 194.310 1831.975 ;
        RECT 5.330 1823.705 194.310 1826.535 ;
        RECT 5.330 1818.265 194.310 1821.095 ;
        RECT 5.330 1812.825 194.310 1815.655 ;
        RECT 5.330 1807.385 194.310 1810.215 ;
        RECT 5.330 1801.945 194.310 1804.775 ;
        RECT 5.330 1796.505 194.310 1799.335 ;
        RECT 5.330 1791.065 194.310 1793.895 ;
        RECT 5.330 1785.625 194.310 1788.455 ;
        RECT 5.330 1780.185 194.310 1783.015 ;
        RECT 5.330 1774.745 194.310 1777.575 ;
        RECT 5.330 1769.305 194.310 1772.135 ;
        RECT 5.330 1763.865 194.310 1766.695 ;
        RECT 5.330 1758.425 194.310 1761.255 ;
        RECT 5.330 1752.985 194.310 1755.815 ;
        RECT 5.330 1747.545 194.310 1750.375 ;
        RECT 5.330 1742.105 194.310 1744.935 ;
        RECT 5.330 1736.665 194.310 1739.495 ;
        RECT 5.330 1731.225 194.310 1734.055 ;
        RECT 5.330 1725.785 194.310 1728.615 ;
        RECT 5.330 1720.345 194.310 1723.175 ;
        RECT 5.330 1714.905 194.310 1717.735 ;
        RECT 5.330 1709.465 194.310 1712.295 ;
        RECT 5.330 1704.025 194.310 1706.855 ;
        RECT 5.330 1698.585 194.310 1701.415 ;
        RECT 5.330 1693.145 194.310 1695.975 ;
        RECT 5.330 1687.705 194.310 1690.535 ;
        RECT 5.330 1682.265 194.310 1685.095 ;
        RECT 5.330 1676.825 194.310 1679.655 ;
        RECT 5.330 1671.385 194.310 1674.215 ;
        RECT 5.330 1665.945 194.310 1668.775 ;
        RECT 5.330 1660.505 194.310 1663.335 ;
        RECT 5.330 1655.065 194.310 1657.895 ;
        RECT 5.330 1649.625 194.310 1652.455 ;
        RECT 5.330 1644.185 194.310 1647.015 ;
        RECT 5.330 1638.745 194.310 1641.575 ;
        RECT 5.330 1633.305 194.310 1636.135 ;
        RECT 5.330 1627.865 194.310 1630.695 ;
        RECT 5.330 1622.425 194.310 1625.255 ;
        RECT 5.330 1616.985 194.310 1619.815 ;
        RECT 5.330 1611.545 194.310 1614.375 ;
        RECT 5.330 1606.105 194.310 1608.935 ;
        RECT 5.330 1600.665 194.310 1603.495 ;
        RECT 5.330 1595.225 194.310 1598.055 ;
        RECT 5.330 1589.785 194.310 1592.615 ;
        RECT 5.330 1584.345 194.310 1587.175 ;
        RECT 5.330 1578.905 194.310 1581.735 ;
        RECT 5.330 1573.465 194.310 1576.295 ;
        RECT 5.330 1568.025 194.310 1570.855 ;
        RECT 5.330 1562.585 194.310 1565.415 ;
        RECT 5.330 1557.145 194.310 1559.975 ;
        RECT 5.330 1551.705 194.310 1554.535 ;
        RECT 5.330 1546.265 194.310 1549.095 ;
        RECT 5.330 1540.825 194.310 1543.655 ;
        RECT 5.330 1535.385 194.310 1538.215 ;
        RECT 5.330 1529.945 194.310 1532.775 ;
        RECT 5.330 1524.505 194.310 1527.335 ;
        RECT 5.330 1519.065 194.310 1521.895 ;
        RECT 5.330 1513.625 194.310 1516.455 ;
        RECT 5.330 1508.185 194.310 1511.015 ;
        RECT 5.330 1502.745 194.310 1505.575 ;
        RECT 5.330 1497.305 194.310 1500.135 ;
        RECT 5.330 1491.865 194.310 1494.695 ;
        RECT 5.330 1486.425 194.310 1489.255 ;
        RECT 5.330 1480.985 194.310 1483.815 ;
        RECT 5.330 1475.545 194.310 1478.375 ;
        RECT 5.330 1470.105 194.310 1472.935 ;
        RECT 5.330 1464.665 194.310 1467.495 ;
        RECT 5.330 1459.225 194.310 1462.055 ;
        RECT 5.330 1453.785 194.310 1456.615 ;
        RECT 5.330 1448.345 194.310 1451.175 ;
        RECT 5.330 1442.905 194.310 1445.735 ;
        RECT 5.330 1437.465 194.310 1440.295 ;
        RECT 5.330 1432.025 194.310 1434.855 ;
        RECT 5.330 1426.585 194.310 1429.415 ;
        RECT 5.330 1421.145 194.310 1423.975 ;
        RECT 5.330 1415.705 194.310 1418.535 ;
        RECT 5.330 1410.265 194.310 1413.095 ;
        RECT 5.330 1404.825 194.310 1407.655 ;
        RECT 5.330 1399.385 194.310 1402.215 ;
        RECT 5.330 1393.945 194.310 1396.775 ;
        RECT 5.330 1388.505 194.310 1391.335 ;
        RECT 5.330 1383.065 194.310 1385.895 ;
        RECT 5.330 1377.625 194.310 1380.455 ;
        RECT 5.330 1372.185 194.310 1375.015 ;
        RECT 5.330 1366.745 194.310 1369.575 ;
        RECT 5.330 1361.305 194.310 1364.135 ;
        RECT 5.330 1355.865 194.310 1358.695 ;
        RECT 5.330 1350.425 194.310 1353.255 ;
        RECT 5.330 1344.985 194.310 1347.815 ;
        RECT 5.330 1339.545 194.310 1342.375 ;
        RECT 5.330 1334.105 194.310 1336.935 ;
        RECT 5.330 1328.665 194.310 1331.495 ;
        RECT 5.330 1323.225 194.310 1326.055 ;
        RECT 5.330 1317.785 194.310 1320.615 ;
        RECT 5.330 1312.345 194.310 1315.175 ;
        RECT 5.330 1306.905 194.310 1309.735 ;
        RECT 5.330 1301.465 194.310 1304.295 ;
        RECT 5.330 1296.025 194.310 1298.855 ;
        RECT 5.330 1290.585 194.310 1293.415 ;
        RECT 5.330 1285.145 194.310 1287.975 ;
        RECT 5.330 1279.705 194.310 1282.535 ;
        RECT 5.330 1274.265 194.310 1277.095 ;
        RECT 5.330 1268.825 194.310 1271.655 ;
        RECT 5.330 1263.385 194.310 1266.215 ;
        RECT 5.330 1257.945 194.310 1260.775 ;
        RECT 5.330 1252.505 194.310 1255.335 ;
        RECT 5.330 1247.065 194.310 1249.895 ;
        RECT 5.330 1241.625 194.310 1244.455 ;
        RECT 5.330 1236.185 194.310 1239.015 ;
        RECT 5.330 1230.745 194.310 1233.575 ;
        RECT 5.330 1225.305 194.310 1228.135 ;
        RECT 5.330 1219.865 194.310 1222.695 ;
        RECT 5.330 1214.425 194.310 1217.255 ;
        RECT 5.330 1208.985 194.310 1211.815 ;
        RECT 5.330 1203.545 194.310 1206.375 ;
        RECT 5.330 1198.105 194.310 1200.935 ;
        RECT 5.330 1192.665 194.310 1195.495 ;
        RECT 5.330 1187.225 194.310 1190.055 ;
        RECT 5.330 1181.785 194.310 1184.615 ;
        RECT 5.330 1176.345 194.310 1179.175 ;
        RECT 5.330 1170.905 194.310 1173.735 ;
        RECT 5.330 1165.465 194.310 1168.295 ;
        RECT 5.330 1160.025 194.310 1162.855 ;
        RECT 5.330 1154.585 194.310 1157.415 ;
        RECT 5.330 1149.145 194.310 1151.975 ;
        RECT 5.330 1143.705 194.310 1146.535 ;
        RECT 5.330 1138.265 194.310 1141.095 ;
        RECT 5.330 1132.825 194.310 1135.655 ;
        RECT 5.330 1127.385 194.310 1130.215 ;
        RECT 5.330 1121.945 194.310 1124.775 ;
        RECT 5.330 1116.505 194.310 1119.335 ;
        RECT 5.330 1111.065 194.310 1113.895 ;
        RECT 5.330 1105.625 194.310 1108.455 ;
        RECT 5.330 1100.185 194.310 1103.015 ;
        RECT 5.330 1094.745 194.310 1097.575 ;
        RECT 5.330 1089.305 194.310 1092.135 ;
        RECT 5.330 1083.865 194.310 1086.695 ;
        RECT 5.330 1078.425 194.310 1081.255 ;
        RECT 5.330 1072.985 194.310 1075.815 ;
        RECT 5.330 1067.545 194.310 1070.375 ;
        RECT 5.330 1062.105 194.310 1064.935 ;
        RECT 5.330 1056.665 194.310 1059.495 ;
        RECT 5.330 1051.225 194.310 1054.055 ;
        RECT 5.330 1045.785 194.310 1048.615 ;
        RECT 5.330 1040.345 194.310 1043.175 ;
        RECT 5.330 1034.905 194.310 1037.735 ;
        RECT 5.330 1029.465 194.310 1032.295 ;
        RECT 5.330 1024.025 194.310 1026.855 ;
        RECT 5.330 1018.585 194.310 1021.415 ;
        RECT 5.330 1013.145 194.310 1015.975 ;
        RECT 5.330 1007.705 194.310 1010.535 ;
        RECT 5.330 1002.265 194.310 1005.095 ;
        RECT 5.330 996.825 194.310 999.655 ;
        RECT 5.330 991.385 194.310 994.215 ;
        RECT 5.330 985.945 194.310 988.775 ;
        RECT 5.330 980.505 194.310 983.335 ;
        RECT 5.330 975.065 194.310 977.895 ;
        RECT 5.330 969.625 194.310 972.455 ;
        RECT 5.330 964.185 194.310 967.015 ;
        RECT 5.330 958.745 194.310 961.575 ;
        RECT 5.330 953.305 194.310 956.135 ;
        RECT 5.330 947.865 194.310 950.695 ;
        RECT 5.330 942.425 194.310 945.255 ;
        RECT 5.330 936.985 194.310 939.815 ;
        RECT 5.330 931.545 194.310 934.375 ;
        RECT 5.330 926.105 194.310 928.935 ;
        RECT 5.330 920.665 194.310 923.495 ;
        RECT 5.330 915.225 194.310 918.055 ;
        RECT 5.330 909.785 194.310 912.615 ;
        RECT 5.330 904.345 194.310 907.175 ;
        RECT 5.330 898.905 194.310 901.735 ;
        RECT 5.330 893.465 194.310 896.295 ;
        RECT 5.330 888.025 194.310 890.855 ;
        RECT 5.330 882.585 194.310 885.415 ;
        RECT 5.330 877.145 194.310 879.975 ;
        RECT 5.330 871.705 194.310 874.535 ;
        RECT 5.330 866.265 194.310 869.095 ;
        RECT 5.330 860.825 194.310 863.655 ;
        RECT 5.330 855.385 194.310 858.215 ;
        RECT 5.330 849.945 194.310 852.775 ;
        RECT 5.330 844.505 194.310 847.335 ;
        RECT 5.330 839.065 194.310 841.895 ;
        RECT 5.330 833.625 194.310 836.455 ;
        RECT 5.330 828.185 194.310 831.015 ;
        RECT 5.330 822.745 194.310 825.575 ;
        RECT 5.330 817.305 194.310 820.135 ;
        RECT 5.330 811.865 194.310 814.695 ;
        RECT 5.330 806.425 194.310 809.255 ;
        RECT 5.330 800.985 194.310 803.815 ;
        RECT 5.330 795.545 194.310 798.375 ;
        RECT 5.330 790.105 194.310 792.935 ;
        RECT 5.330 784.665 194.310 787.495 ;
        RECT 5.330 779.225 194.310 782.055 ;
        RECT 5.330 773.785 194.310 776.615 ;
        RECT 5.330 768.345 194.310 771.175 ;
        RECT 5.330 762.905 194.310 765.735 ;
        RECT 5.330 757.465 194.310 760.295 ;
        RECT 5.330 752.025 194.310 754.855 ;
        RECT 5.330 746.585 194.310 749.415 ;
        RECT 5.330 741.145 194.310 743.975 ;
        RECT 5.330 735.705 194.310 738.535 ;
        RECT 5.330 730.265 194.310 733.095 ;
        RECT 5.330 724.825 194.310 727.655 ;
        RECT 5.330 719.385 194.310 722.215 ;
        RECT 5.330 713.945 194.310 716.775 ;
        RECT 5.330 708.505 194.310 711.335 ;
        RECT 5.330 703.065 194.310 705.895 ;
        RECT 5.330 697.625 194.310 700.455 ;
        RECT 5.330 692.185 194.310 695.015 ;
        RECT 5.330 686.745 194.310 689.575 ;
        RECT 5.330 681.305 194.310 684.135 ;
        RECT 5.330 675.865 194.310 678.695 ;
        RECT 5.330 670.425 194.310 673.255 ;
        RECT 5.330 664.985 194.310 667.815 ;
        RECT 5.330 659.545 194.310 662.375 ;
        RECT 5.330 654.105 194.310 656.935 ;
        RECT 5.330 648.665 194.310 651.495 ;
        RECT 5.330 643.225 194.310 646.055 ;
        RECT 5.330 637.785 194.310 640.615 ;
        RECT 5.330 632.345 194.310 635.175 ;
        RECT 5.330 626.905 194.310 629.735 ;
        RECT 5.330 621.465 194.310 624.295 ;
        RECT 5.330 616.025 194.310 618.855 ;
        RECT 5.330 610.585 194.310 613.415 ;
        RECT 5.330 605.145 194.310 607.975 ;
        RECT 5.330 599.705 194.310 602.535 ;
        RECT 5.330 594.265 194.310 597.095 ;
        RECT 5.330 588.825 194.310 591.655 ;
        RECT 5.330 583.385 194.310 586.215 ;
        RECT 5.330 577.945 194.310 580.775 ;
        RECT 5.330 572.505 194.310 575.335 ;
        RECT 5.330 567.065 194.310 569.895 ;
        RECT 5.330 561.625 194.310 564.455 ;
        RECT 5.330 556.185 194.310 559.015 ;
        RECT 5.330 550.745 194.310 553.575 ;
        RECT 5.330 545.305 194.310 548.135 ;
        RECT 5.330 539.865 194.310 542.695 ;
        RECT 5.330 534.425 194.310 537.255 ;
        RECT 5.330 528.985 194.310 531.815 ;
        RECT 5.330 523.545 194.310 526.375 ;
        RECT 5.330 518.105 194.310 520.935 ;
        RECT 5.330 512.665 194.310 515.495 ;
        RECT 5.330 507.225 194.310 510.055 ;
        RECT 5.330 501.785 194.310 504.615 ;
        RECT 5.330 496.345 194.310 499.175 ;
        RECT 5.330 490.905 194.310 493.735 ;
        RECT 5.330 485.465 194.310 488.295 ;
        RECT 5.330 480.025 194.310 482.855 ;
        RECT 5.330 474.585 194.310 477.415 ;
        RECT 5.330 469.145 194.310 471.975 ;
        RECT 5.330 463.705 194.310 466.535 ;
        RECT 5.330 458.265 194.310 461.095 ;
        RECT 5.330 452.825 194.310 455.655 ;
        RECT 5.330 447.385 194.310 450.215 ;
        RECT 5.330 441.945 194.310 444.775 ;
        RECT 5.330 436.505 194.310 439.335 ;
        RECT 5.330 431.065 194.310 433.895 ;
        RECT 5.330 425.625 194.310 428.455 ;
        RECT 5.330 420.185 194.310 423.015 ;
        RECT 5.330 414.745 194.310 417.575 ;
        RECT 5.330 409.305 194.310 412.135 ;
        RECT 5.330 403.865 194.310 406.695 ;
        RECT 5.330 398.425 194.310 401.255 ;
        RECT 5.330 392.985 194.310 395.815 ;
        RECT 5.330 387.545 194.310 390.375 ;
        RECT 5.330 382.105 194.310 384.935 ;
        RECT 5.330 376.665 194.310 379.495 ;
        RECT 5.330 371.225 194.310 374.055 ;
        RECT 5.330 365.785 194.310 368.615 ;
        RECT 5.330 360.345 194.310 363.175 ;
        RECT 5.330 354.905 194.310 357.735 ;
        RECT 5.330 349.465 194.310 352.295 ;
        RECT 5.330 344.025 194.310 346.855 ;
        RECT 5.330 338.585 194.310 341.415 ;
        RECT 5.330 333.145 194.310 335.975 ;
        RECT 5.330 327.705 194.310 330.535 ;
        RECT 5.330 322.265 194.310 325.095 ;
        RECT 5.330 316.825 194.310 319.655 ;
        RECT 5.330 311.385 194.310 314.215 ;
        RECT 5.330 305.945 194.310 308.775 ;
        RECT 5.330 300.505 194.310 303.335 ;
        RECT 5.330 295.065 194.310 297.895 ;
        RECT 5.330 289.625 194.310 292.455 ;
        RECT 5.330 284.185 194.310 287.015 ;
        RECT 5.330 278.745 194.310 281.575 ;
        RECT 5.330 273.305 194.310 276.135 ;
        RECT 5.330 267.865 194.310 270.695 ;
        RECT 5.330 262.425 194.310 265.255 ;
        RECT 5.330 256.985 194.310 259.815 ;
        RECT 5.330 251.545 194.310 254.375 ;
        RECT 5.330 246.105 194.310 248.935 ;
        RECT 5.330 240.665 194.310 243.495 ;
        RECT 5.330 235.225 194.310 238.055 ;
        RECT 5.330 229.785 194.310 232.615 ;
        RECT 5.330 224.345 194.310 227.175 ;
        RECT 5.330 218.905 194.310 221.735 ;
        RECT 5.330 213.465 194.310 216.295 ;
        RECT 5.330 208.025 194.310 210.855 ;
        RECT 5.330 202.585 194.310 205.415 ;
        RECT 5.330 197.145 194.310 199.975 ;
        RECT 5.330 191.705 194.310 194.535 ;
        RECT 5.330 186.265 194.310 189.095 ;
        RECT 5.330 180.825 194.310 183.655 ;
        RECT 5.330 175.385 194.310 178.215 ;
        RECT 5.330 169.945 194.310 172.775 ;
        RECT 5.330 164.505 194.310 167.335 ;
        RECT 5.330 159.065 194.310 161.895 ;
        RECT 5.330 153.625 194.310 156.455 ;
        RECT 5.330 148.185 194.310 151.015 ;
        RECT 5.330 142.745 194.310 145.575 ;
        RECT 5.330 137.305 194.310 140.135 ;
        RECT 5.330 131.865 194.310 134.695 ;
        RECT 5.330 126.425 194.310 129.255 ;
        RECT 5.330 120.985 194.310 123.815 ;
        RECT 5.330 115.545 194.310 118.375 ;
        RECT 5.330 110.105 194.310 112.935 ;
        RECT 5.330 104.665 194.310 107.495 ;
        RECT 5.330 99.225 194.310 102.055 ;
        RECT 5.330 93.785 194.310 96.615 ;
        RECT 5.330 88.345 194.310 91.175 ;
        RECT 5.330 82.905 194.310 85.735 ;
        RECT 5.330 77.465 194.310 80.295 ;
        RECT 5.330 72.025 194.310 74.855 ;
        RECT 5.330 66.585 194.310 69.415 ;
        RECT 5.330 61.145 194.310 63.975 ;
        RECT 5.330 55.705 194.310 58.535 ;
        RECT 5.330 50.265 194.310 53.095 ;
        RECT 5.330 44.825 194.310 47.655 ;
        RECT 5.330 39.385 194.310 42.215 ;
        RECT 5.330 33.945 194.310 36.775 ;
        RECT 5.330 28.505 194.310 31.335 ;
        RECT 5.330 23.065 194.310 25.895 ;
        RECT 5.330 17.625 194.310 20.455 ;
        RECT 5.330 12.185 194.310 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 194.120 2986.645 ;
      LAYER met1 ;
        RECT 5.520 10.640 194.120 2986.800 ;
      LAYER met2 ;
        RECT 21.070 4.280 192.650 2986.745 ;
        RECT 21.070 4.000 49.490 4.280 ;
        RECT 50.330 4.000 149.310 4.280 ;
        RECT 150.150 4.000 192.650 4.280 ;
      LAYER met3 ;
        RECT 21.050 2899.200 196.000 2986.725 ;
        RECT 21.050 2897.800 195.600 2899.200 ;
        RECT 21.050 2699.280 196.000 2897.800 ;
        RECT 21.050 2697.880 195.600 2699.280 ;
        RECT 21.050 2499.360 196.000 2697.880 ;
        RECT 21.050 2497.960 195.600 2499.360 ;
        RECT 21.050 2299.440 196.000 2497.960 ;
        RECT 21.050 2298.040 195.600 2299.440 ;
        RECT 21.050 2099.520 196.000 2298.040 ;
        RECT 21.050 2098.120 195.600 2099.520 ;
        RECT 21.050 1899.600 196.000 2098.120 ;
        RECT 21.050 1898.200 195.600 1899.600 ;
        RECT 21.050 1699.680 196.000 1898.200 ;
        RECT 21.050 1698.280 195.600 1699.680 ;
        RECT 21.050 1499.760 196.000 1698.280 ;
        RECT 21.050 1498.360 195.600 1499.760 ;
        RECT 21.050 1299.840 196.000 1498.360 ;
        RECT 21.050 1298.440 195.600 1299.840 ;
        RECT 21.050 1099.920 196.000 1298.440 ;
        RECT 21.050 1098.520 195.600 1099.920 ;
        RECT 21.050 900.000 196.000 1098.520 ;
        RECT 21.050 898.600 195.600 900.000 ;
        RECT 21.050 700.080 196.000 898.600 ;
        RECT 21.050 698.680 195.600 700.080 ;
        RECT 21.050 500.160 196.000 698.680 ;
        RECT 21.050 498.760 195.600 500.160 ;
        RECT 21.050 300.240 196.000 498.760 ;
        RECT 21.050 298.840 195.600 300.240 ;
        RECT 21.050 100.320 196.000 298.840 ;
        RECT 21.050 98.920 195.600 100.320 ;
        RECT 21.050 10.715 196.000 98.920 ;
  END
END user_proj_example
END LIBRARY

