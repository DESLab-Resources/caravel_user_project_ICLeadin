magic
tech sky130A
magscale 1 2
timestamp 1727667461
<< nwell >>
rect 1066 596485 38862 597051
rect 1066 595397 38862 595963
rect 1066 594309 38862 594875
rect 1066 593221 38862 593787
rect 1066 592133 38862 592699
rect 1066 591045 38862 591611
rect 1066 589957 38862 590523
rect 1066 588869 38862 589435
rect 1066 587781 38862 588347
rect 1066 586693 38862 587259
rect 1066 585605 38862 586171
rect 1066 584517 38862 585083
rect 1066 583429 38862 583995
rect 1066 582341 38862 582907
rect 1066 581253 38862 581819
rect 1066 580165 38862 580731
rect 1066 579077 38862 579643
rect 1066 577989 38862 578555
rect 1066 576901 38862 577467
rect 1066 575813 38862 576379
rect 1066 574725 38862 575291
rect 1066 573637 38862 574203
rect 1066 572549 38862 573115
rect 1066 571461 38862 572027
rect 1066 570373 38862 570939
rect 1066 569285 38862 569851
rect 1066 568197 38862 568763
rect 1066 567109 38862 567675
rect 1066 566021 38862 566587
rect 1066 564933 38862 565499
rect 1066 563845 38862 564411
rect 1066 562757 38862 563323
rect 1066 561669 38862 562235
rect 1066 560581 38862 561147
rect 1066 559493 38862 560059
rect 1066 558405 38862 558971
rect 1066 557317 38862 557883
rect 1066 556229 38862 556795
rect 1066 555141 38862 555707
rect 1066 554053 38862 554619
rect 1066 552965 38862 553531
rect 1066 551877 38862 552443
rect 1066 550789 38862 551355
rect 1066 549701 38862 550267
rect 1066 548613 38862 549179
rect 1066 547525 38862 548091
rect 1066 546437 38862 547003
rect 1066 545349 38862 545915
rect 1066 544261 38862 544827
rect 1066 543173 38862 543739
rect 1066 542085 38862 542651
rect 1066 540997 38862 541563
rect 1066 539909 38862 540475
rect 1066 538821 38862 539387
rect 1066 537733 38862 538299
rect 1066 536645 38862 537211
rect 1066 535557 38862 536123
rect 1066 534469 38862 535035
rect 1066 533381 38862 533947
rect 1066 532293 38862 532859
rect 1066 531205 38862 531771
rect 1066 530117 38862 530683
rect 1066 529029 38862 529595
rect 1066 527941 38862 528507
rect 1066 526853 38862 527419
rect 1066 525765 38862 526331
rect 1066 524677 38862 525243
rect 1066 523589 38862 524155
rect 1066 522501 38862 523067
rect 1066 521413 38862 521979
rect 1066 520325 38862 520891
rect 1066 519237 38862 519803
rect 1066 518149 38862 518715
rect 1066 517061 38862 517627
rect 1066 515973 38862 516539
rect 1066 514885 38862 515451
rect 1066 513797 38862 514363
rect 1066 512709 38862 513275
rect 1066 511621 38862 512187
rect 1066 510533 38862 511099
rect 1066 509445 38862 510011
rect 1066 508357 38862 508923
rect 1066 507269 38862 507835
rect 1066 506181 38862 506747
rect 1066 505093 38862 505659
rect 1066 504005 38862 504571
rect 1066 502917 38862 503483
rect 1066 501829 38862 502395
rect 1066 500741 38862 501307
rect 1066 499653 38862 500219
rect 1066 498565 38862 499131
rect 1066 497477 38862 498043
rect 1066 496389 38862 496955
rect 1066 495301 38862 495867
rect 1066 494213 38862 494779
rect 1066 493125 38862 493691
rect 1066 492037 38862 492603
rect 1066 490949 38862 491515
rect 1066 489861 38862 490427
rect 1066 488773 38862 489339
rect 1066 487685 38862 488251
rect 1066 486597 38862 487163
rect 1066 485509 38862 486075
rect 1066 484421 38862 484987
rect 1066 483333 38862 483899
rect 1066 482245 38862 482811
rect 1066 481157 38862 481723
rect 1066 480069 38862 480635
rect 1066 478981 38862 479547
rect 1066 477893 38862 478459
rect 1066 476805 38862 477371
rect 1066 475717 38862 476283
rect 1066 474629 38862 475195
rect 1066 473541 38862 474107
rect 1066 472453 38862 473019
rect 1066 471365 38862 471931
rect 1066 470277 38862 470843
rect 1066 469189 38862 469755
rect 1066 468101 38862 468667
rect 1066 467013 38862 467579
rect 1066 465925 38862 466491
rect 1066 464837 38862 465403
rect 1066 463749 38862 464315
rect 1066 462661 38862 463227
rect 1066 461573 38862 462139
rect 1066 460485 38862 461051
rect 1066 459397 38862 459963
rect 1066 458309 38862 458875
rect 1066 457221 38862 457787
rect 1066 456133 38862 456699
rect 1066 455045 38862 455611
rect 1066 453957 38862 454523
rect 1066 452869 38862 453435
rect 1066 451781 38862 452347
rect 1066 450693 38862 451259
rect 1066 449605 38862 450171
rect 1066 448517 38862 449083
rect 1066 447429 38862 447995
rect 1066 446341 38862 446907
rect 1066 445253 38862 445819
rect 1066 444165 38862 444731
rect 1066 443077 38862 443643
rect 1066 441989 38862 442555
rect 1066 440901 38862 441467
rect 1066 439813 38862 440379
rect 1066 438725 38862 439291
rect 1066 437637 38862 438203
rect 1066 436549 38862 437115
rect 1066 435461 38862 436027
rect 1066 434373 38862 434939
rect 1066 433285 38862 433851
rect 1066 432197 38862 432763
rect 1066 431109 38862 431675
rect 1066 430021 38862 430587
rect 1066 428933 38862 429499
rect 1066 427845 38862 428411
rect 1066 426757 38862 427323
rect 1066 425669 38862 426235
rect 1066 424581 38862 425147
rect 1066 423493 38862 424059
rect 1066 422405 38862 422971
rect 1066 421317 38862 421883
rect 1066 420229 38862 420795
rect 1066 419141 38862 419707
rect 1066 418053 38862 418619
rect 1066 416965 38862 417531
rect 1066 415877 38862 416443
rect 1066 414789 38862 415355
rect 1066 413701 38862 414267
rect 1066 412613 38862 413179
rect 1066 411525 38862 412091
rect 1066 410437 38862 411003
rect 1066 409349 38862 409915
rect 1066 408261 38862 408827
rect 1066 407173 38862 407739
rect 1066 406085 38862 406651
rect 1066 404997 38862 405563
rect 1066 403909 38862 404475
rect 1066 402821 38862 403387
rect 1066 401733 38862 402299
rect 1066 400645 38862 401211
rect 1066 399557 38862 400123
rect 1066 398469 38862 399035
rect 1066 397381 38862 397947
rect 1066 396293 38862 396859
rect 1066 395205 38862 395771
rect 1066 394117 38862 394683
rect 1066 393029 38862 393595
rect 1066 391941 38862 392507
rect 1066 390853 38862 391419
rect 1066 389765 38862 390331
rect 1066 388677 38862 389243
rect 1066 387589 38862 388155
rect 1066 386501 38862 387067
rect 1066 385413 38862 385979
rect 1066 384325 38862 384891
rect 1066 383237 38862 383803
rect 1066 382149 38862 382715
rect 1066 381061 38862 381627
rect 1066 379973 38862 380539
rect 1066 378885 38862 379451
rect 1066 377797 38862 378363
rect 1066 376709 38862 377275
rect 1066 375621 38862 376187
rect 1066 374533 38862 375099
rect 1066 373445 38862 374011
rect 1066 372357 38862 372923
rect 1066 371269 38862 371835
rect 1066 370181 38862 370747
rect 1066 369093 38862 369659
rect 1066 368005 38862 368571
rect 1066 366917 38862 367483
rect 1066 365829 38862 366395
rect 1066 364741 38862 365307
rect 1066 363653 38862 364219
rect 1066 362565 38862 363131
rect 1066 361477 38862 362043
rect 1066 360389 38862 360955
rect 1066 359301 38862 359867
rect 1066 358213 38862 358779
rect 1066 357125 38862 357691
rect 1066 356037 38862 356603
rect 1066 354949 38862 355515
rect 1066 353861 38862 354427
rect 1066 352773 38862 353339
rect 1066 351685 38862 352251
rect 1066 350597 38862 351163
rect 1066 349509 38862 350075
rect 1066 348421 38862 348987
rect 1066 347333 38862 347899
rect 1066 346245 38862 346811
rect 1066 345157 38862 345723
rect 1066 344069 38862 344635
rect 1066 342981 38862 343547
rect 1066 341893 38862 342459
rect 1066 340805 38862 341371
rect 1066 339717 38862 340283
rect 1066 338629 38862 339195
rect 1066 337541 38862 338107
rect 1066 336453 38862 337019
rect 1066 335365 38862 335931
rect 1066 334277 38862 334843
rect 1066 333189 38862 333755
rect 1066 332101 38862 332667
rect 1066 331013 38862 331579
rect 1066 329925 38862 330491
rect 1066 328837 38862 329403
rect 1066 327749 38862 328315
rect 1066 326661 38862 327227
rect 1066 325573 38862 326139
rect 1066 324485 38862 325051
rect 1066 323397 38862 323963
rect 1066 322309 38862 322875
rect 1066 321221 38862 321787
rect 1066 320133 38862 320699
rect 1066 319045 38862 319611
rect 1066 317957 38862 318523
rect 1066 316869 38862 317435
rect 1066 315781 38862 316347
rect 1066 314693 38862 315259
rect 1066 313605 38862 314171
rect 1066 312517 38862 313083
rect 1066 311429 38862 311995
rect 1066 310341 38862 310907
rect 1066 309253 38862 309819
rect 1066 308165 38862 308731
rect 1066 307077 38862 307643
rect 1066 305989 38862 306555
rect 1066 304901 38862 305467
rect 1066 303813 38862 304379
rect 1066 302725 38862 303291
rect 1066 301637 38862 302203
rect 1066 300549 38862 301115
rect 1066 299461 38862 300027
rect 1066 298373 38862 298939
rect 1066 297285 38862 297851
rect 1066 296197 38862 296763
rect 1066 295109 38862 295675
rect 1066 294021 38862 294587
rect 1066 292933 38862 293499
rect 1066 291845 38862 292411
rect 1066 290757 38862 291323
rect 1066 289669 38862 290235
rect 1066 288581 38862 289147
rect 1066 287493 38862 288059
rect 1066 286405 38862 286971
rect 1066 285317 38862 285883
rect 1066 284229 38862 284795
rect 1066 283141 38862 283707
rect 1066 282053 38862 282619
rect 1066 280965 38862 281531
rect 1066 279877 38862 280443
rect 1066 278789 38862 279355
rect 1066 277701 38862 278267
rect 1066 276613 38862 277179
rect 1066 275525 38862 276091
rect 1066 274437 38862 275003
rect 1066 273349 38862 273915
rect 1066 272261 38862 272827
rect 1066 271173 38862 271739
rect 1066 270085 38862 270651
rect 1066 268997 38862 269563
rect 1066 267909 38862 268475
rect 1066 266821 38862 267387
rect 1066 265733 38862 266299
rect 1066 264645 38862 265211
rect 1066 263557 38862 264123
rect 1066 262469 38862 263035
rect 1066 261381 38862 261947
rect 1066 260293 38862 260859
rect 1066 259205 38862 259771
rect 1066 258117 38862 258683
rect 1066 257029 38862 257595
rect 1066 255941 38862 256507
rect 1066 254853 38862 255419
rect 1066 253765 38862 254331
rect 1066 252677 38862 253243
rect 1066 251589 38862 252155
rect 1066 250501 38862 251067
rect 1066 249413 38862 249979
rect 1066 248325 38862 248891
rect 1066 247237 38862 247803
rect 1066 246149 38862 246715
rect 1066 245061 38862 245627
rect 1066 243973 38862 244539
rect 1066 242885 38862 243451
rect 1066 241797 38862 242363
rect 1066 240709 38862 241275
rect 1066 239621 38862 240187
rect 1066 238533 38862 239099
rect 1066 237445 38862 238011
rect 1066 236357 38862 236923
rect 1066 235269 38862 235835
rect 1066 234181 38862 234747
rect 1066 233093 38862 233659
rect 1066 232005 38862 232571
rect 1066 230917 38862 231483
rect 1066 229829 38862 230395
rect 1066 228741 38862 229307
rect 1066 227653 38862 228219
rect 1066 226565 38862 227131
rect 1066 225477 38862 226043
rect 1066 224389 38862 224955
rect 1066 223301 38862 223867
rect 1066 222213 38862 222779
rect 1066 221125 38862 221691
rect 1066 220037 38862 220603
rect 1066 218949 38862 219515
rect 1066 217861 38862 218427
rect 1066 216773 38862 217339
rect 1066 215685 38862 216251
rect 1066 214597 38862 215163
rect 1066 213509 38862 214075
rect 1066 212421 38862 212987
rect 1066 211333 38862 211899
rect 1066 210245 38862 210811
rect 1066 209157 38862 209723
rect 1066 208069 38862 208635
rect 1066 206981 38862 207547
rect 1066 205893 38862 206459
rect 1066 204805 38862 205371
rect 1066 203717 38862 204283
rect 1066 202629 38862 203195
rect 1066 201541 38862 202107
rect 1066 200453 38862 201019
rect 1066 199365 38862 199931
rect 1066 198277 38862 198843
rect 1066 197189 38862 197755
rect 1066 196101 38862 196667
rect 1066 195013 38862 195579
rect 1066 193925 38862 194491
rect 1066 192837 38862 193403
rect 1066 191749 38862 192315
rect 1066 190661 38862 191227
rect 1066 189573 38862 190139
rect 1066 188485 38862 189051
rect 1066 187397 38862 187963
rect 1066 186309 38862 186875
rect 1066 185221 38862 185787
rect 1066 184133 38862 184699
rect 1066 183045 38862 183611
rect 1066 181957 38862 182523
rect 1066 180869 38862 181435
rect 1066 179781 38862 180347
rect 1066 178693 38862 179259
rect 1066 177605 38862 178171
rect 1066 176517 38862 177083
rect 1066 175429 38862 175995
rect 1066 174341 38862 174907
rect 1066 173253 38862 173819
rect 1066 172165 38862 172731
rect 1066 171077 38862 171643
rect 1066 169989 38862 170555
rect 1066 168901 38862 169467
rect 1066 167813 38862 168379
rect 1066 166725 38862 167291
rect 1066 165637 38862 166203
rect 1066 164549 38862 165115
rect 1066 163461 38862 164027
rect 1066 162373 38862 162939
rect 1066 161285 38862 161851
rect 1066 160197 38862 160763
rect 1066 159109 38862 159675
rect 1066 158021 38862 158587
rect 1066 156933 38862 157499
rect 1066 155845 38862 156411
rect 1066 154757 38862 155323
rect 1066 153669 38862 154235
rect 1066 152581 38862 153147
rect 1066 151493 38862 152059
rect 1066 150405 38862 150971
rect 1066 149317 38862 149883
rect 1066 148229 38862 148795
rect 1066 147141 38862 147707
rect 1066 146053 38862 146619
rect 1066 144965 38862 145531
rect 1066 143877 38862 144443
rect 1066 142789 38862 143355
rect 1066 141701 38862 142267
rect 1066 140613 38862 141179
rect 1066 139525 38862 140091
rect 1066 138437 38862 139003
rect 1066 137349 38862 137915
rect 1066 136261 38862 136827
rect 1066 135173 38862 135739
rect 1066 134085 38862 134651
rect 1066 132997 38862 133563
rect 1066 131909 38862 132475
rect 1066 130821 38862 131387
rect 1066 129733 38862 130299
rect 1066 128645 38862 129211
rect 1066 127557 38862 128123
rect 1066 126469 38862 127035
rect 1066 125381 38862 125947
rect 1066 124293 38862 124859
rect 1066 123205 38862 123771
rect 1066 122117 38862 122683
rect 1066 121029 38862 121595
rect 1066 119941 38862 120507
rect 1066 118853 38862 119419
rect 1066 117765 38862 118331
rect 1066 116677 38862 117243
rect 1066 115589 38862 116155
rect 1066 114501 38862 115067
rect 1066 113413 38862 113979
rect 1066 112325 38862 112891
rect 1066 111237 38862 111803
rect 1066 110149 38862 110715
rect 1066 109061 38862 109627
rect 1066 107973 38862 108539
rect 1066 106885 38862 107451
rect 1066 105797 38862 106363
rect 1066 104709 38862 105275
rect 1066 103621 38862 104187
rect 1066 102533 38862 103099
rect 1066 101445 38862 102011
rect 1066 100357 38862 100923
rect 1066 99269 38862 99835
rect 1066 98181 38862 98747
rect 1066 97093 38862 97659
rect 1066 96005 38862 96571
rect 1066 94917 38862 95483
rect 1066 93829 38862 94395
rect 1066 92741 38862 93307
rect 1066 91653 38862 92219
rect 1066 90565 38862 91131
rect 1066 89477 38862 90043
rect 1066 88389 38862 88955
rect 1066 87301 38862 87867
rect 1066 86213 38862 86779
rect 1066 85125 38862 85691
rect 1066 84037 38862 84603
rect 1066 82949 38862 83515
rect 1066 81861 38862 82427
rect 1066 80773 38862 81339
rect 1066 79685 38862 80251
rect 1066 78597 38862 79163
rect 1066 77509 38862 78075
rect 1066 76421 38862 76987
rect 1066 75333 38862 75899
rect 1066 74245 38862 74811
rect 1066 73157 38862 73723
rect 1066 72069 38862 72635
rect 1066 70981 38862 71547
rect 1066 69893 38862 70459
rect 1066 68805 38862 69371
rect 1066 67717 38862 68283
rect 1066 66629 38862 67195
rect 1066 65541 38862 66107
rect 1066 64453 38862 65019
rect 1066 63365 38862 63931
rect 1066 62277 38862 62843
rect 1066 61189 38862 61755
rect 1066 60101 38862 60667
rect 1066 59013 38862 59579
rect 1066 57925 38862 58491
rect 1066 56837 38862 57403
rect 1066 55749 38862 56315
rect 1066 54661 38862 55227
rect 1066 53573 38862 54139
rect 1066 52485 38862 53051
rect 1066 51397 38862 51963
rect 1066 50309 38862 50875
rect 1066 49221 38862 49787
rect 1066 48133 38862 48699
rect 1066 47045 38862 47611
rect 1066 45957 38862 46523
rect 1066 44869 38862 45435
rect 1066 43781 38862 44347
rect 1066 42693 38862 43259
rect 1066 41605 38862 42171
rect 1066 40517 38862 41083
rect 1066 39429 38862 39995
rect 1066 38341 38862 38907
rect 1066 37253 38862 37819
rect 1066 36165 38862 36731
rect 1066 35077 38862 35643
rect 1066 33989 38862 34555
rect 1066 32901 38862 33467
rect 1066 31813 38862 32379
rect 1066 30725 38862 31291
rect 1066 29637 38862 30203
rect 1066 28549 38862 29115
rect 1066 27461 38862 28027
rect 1066 26373 38862 26939
rect 1066 25285 38862 25851
rect 1066 24197 38862 24763
rect 1066 23109 38862 23675
rect 1066 22021 38862 22587
rect 1066 20933 38862 21499
rect 1066 19845 38862 20411
rect 1066 18757 38862 19323
rect 1066 17669 38862 18235
rect 1066 16581 38862 17147
rect 1066 15493 38862 16059
rect 1066 14405 38862 14971
rect 1066 13317 38862 13883
rect 1066 12229 38862 12795
rect 1066 11141 38862 11707
rect 1066 10053 38862 10619
rect 1066 8965 38862 9531
rect 1066 7877 38862 8443
rect 1066 6789 38862 7355
rect 1066 5701 38862 6267
rect 1066 4613 38862 5179
rect 1066 3525 38862 4091
rect 1066 2437 38862 3003
<< obsli1 >>
rect 1104 2159 38824 597329
<< obsm1 >>
rect 1104 2128 38824 597360
<< metal2 >>
rect 9954 0 10010 800
rect 29918 0 29974 800
<< obsm2 >>
rect 4214 856 38530 597349
rect 4214 800 9898 856
rect 10066 800 29862 856
rect 30030 800 38530 856
<< metal3 >>
rect 39200 579640 40000 579760
rect 39200 539656 40000 539776
rect 39200 499672 40000 499792
rect 39200 459688 40000 459808
rect 39200 419704 40000 419824
rect 39200 379720 40000 379840
rect 39200 339736 40000 339856
rect 39200 299752 40000 299872
rect 39200 259768 40000 259888
rect 39200 219784 40000 219904
rect 39200 179800 40000 179920
rect 39200 139816 40000 139936
rect 39200 99832 40000 99952
rect 39200 59848 40000 59968
rect 39200 19864 40000 19984
<< obsm3 >>
rect 4210 579840 39200 597345
rect 4210 579560 39120 579840
rect 4210 539856 39200 579560
rect 4210 539576 39120 539856
rect 4210 499872 39200 539576
rect 4210 499592 39120 499872
rect 4210 459888 39200 499592
rect 4210 459608 39120 459888
rect 4210 419904 39200 459608
rect 4210 419624 39120 419904
rect 4210 379920 39200 419624
rect 4210 379640 39120 379920
rect 4210 339936 39200 379640
rect 4210 339656 39120 339936
rect 4210 299952 39200 339656
rect 4210 299672 39120 299952
rect 4210 259968 39200 299672
rect 4210 259688 39120 259968
rect 4210 219984 39200 259688
rect 4210 219704 39120 219984
rect 4210 180000 39200 219704
rect 4210 179720 39120 180000
rect 4210 140016 39200 179720
rect 4210 139736 39120 140016
rect 4210 100032 39200 139736
rect 4210 99752 39120 100032
rect 4210 60048 39200 99752
rect 4210 59768 39120 60048
rect 4210 20064 39200 59768
rect 4210 19784 39120 20064
rect 4210 2143 39200 19784
<< metal4 >>
rect 4208 2128 4528 597360
rect 19568 2128 19888 597360
rect 34928 2128 35248 597360
<< labels >>
rlabel metal3 s 39200 19864 40000 19984 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 39200 139816 40000 139936 6 io_in[1]
port 2 nsew signal input
rlabel metal3 s 39200 259768 40000 259888 6 io_in[2]
port 3 nsew signal input
rlabel metal3 s 39200 379720 40000 379840 6 io_in[3]
port 4 nsew signal input
rlabel metal3 s 39200 499672 40000 499792 6 io_in[4]
port 5 nsew signal input
rlabel metal3 s 39200 99832 40000 99952 6 io_oeb[0]
port 6 nsew signal output
rlabel metal3 s 39200 219784 40000 219904 6 io_oeb[1]
port 7 nsew signal output
rlabel metal3 s 39200 339736 40000 339856 6 io_oeb[2]
port 8 nsew signal output
rlabel metal3 s 39200 459688 40000 459808 6 io_oeb[3]
port 9 nsew signal output
rlabel metal3 s 39200 579640 40000 579760 6 io_oeb[4]
port 10 nsew signal output
rlabel metal3 s 39200 59848 40000 59968 6 io_out[0]
port 11 nsew signal output
rlabel metal3 s 39200 179800 40000 179920 6 io_out[1]
port 12 nsew signal output
rlabel metal3 s 39200 299752 40000 299872 6 io_out[2]
port 13 nsew signal output
rlabel metal3 s 39200 419704 40000 419824 6 io_out[3]
port 14 nsew signal output
rlabel metal3 s 39200 539656 40000 539776 6 io_out[4]
port 15 nsew signal output
rlabel metal4 s 4208 2128 4528 597360 6 vccd1
port 16 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 597360 6 vccd1
port 16 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 597360 6 vssd1
port 17 nsew ground bidirectional
rlabel metal2 s 9954 0 10010 800 6 wb_clk_i
port 18 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 wb_rst_i
port 19 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 40000 600000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 6481520
string GDS_FILE /home/icuser/caravel_user_project_ICLeadin/openlane/user_proj_example/runs/24_09_30_10_36/results/signoff/user_proj_example.magic.gds
string GDS_START 130200
<< end >>

